//Q74. How can all assertions be turned off during simulation?

NOTE: Same as Question No- 37 , Please refer the answer.
