//Q60. What is a sequence repetition operator? What are the three different type of repetition operators used in sequences in SVA?

In SystemVerilog Assertions (SVA), sequence repetition operators are used to specify how many times a particular event or condition should occur within a sequence.
These operators allow you to define complex temporal behaviors by repeating certain parts of a sequence a specified number of times. 
There are three different types of repetition operators used in sequences in SVA:
   
  1. Consecutive Repetition ([*n ])
  2. Non-Consecutive Repetition ([=n])
  3. Goto Repetition ([->n])
