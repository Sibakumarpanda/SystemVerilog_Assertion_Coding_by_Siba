//Q68. Write an assertion checker to make sure that an output signal never goes X?

NOTE: The solution is same as ( Question No : 9,32,68)
