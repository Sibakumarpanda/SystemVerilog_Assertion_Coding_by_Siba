/*Q65 Are following assertions equivalent?
 a) @(posedge clk) req |=> ##10 $rose(ack);
 b) @(posedge clk) req |-> ##11 $rose(ack); 
 */

Refer Question No 26 and its Solution for this (NOTE: Question No 26 and Question No 65 , both are same)
