//3. Sequence samples values of a and b on every positive edge of clk and evaluates to true if both a and b are equal
module concurrent_example; 
  bit clk;
  bit a,b;
always #5 clk = ~clk; 
initial begin
      a=0; b=0;
  #15 a=1; b=0; //15
  #10 a=0; b=1; //25
  #10 a=0; b=1; //35
  #10 a=0; b=0; //45
  #10 a=0; b=1; //55
  #10 a=0; b=0; //65
  #10 a=0; b=0; //75
  #10 a=1; b=0; //85
  #10 a=0; b=1; //95
  #10 a=0; b=0; //105
  #10 a=0; b=1; //115
  #10 a=0; b=0; //125
  #10 a=0; b=1; //135
  #10 a=0; b=0; //145
  #10 a=0; b=0; //155
  #10;
  $finish;
end

property check_a_b_equal;
  @(posedge clk) 
  (a == b);
endproperty
  
P1:assert property (check_a_b_equal)   
   $display("PASSED at TIME=%0d with a=%0b b= %0b ",$time ,a,b);    
  else      
    $error("FAILED at TIME=%0d with a=%0b b= %0b ",$time ,a,b);

initial begin
   $dumpfile("waveform.vcd");
   $dumpvars();
  end  
  endmodule
  
// Log File output  
[2025-05-04 09:21:01 UTC] vcs -full64 -licqueue '-timescale=1ns/1ns' '+vcs+flush+all' '+warn=all' '-sverilog' design.sv testbench.sv  && ./simv +vcs+lic+wait  
                         Chronologic VCS (TM)
       Version U-2023.03-SP2_Full64 -- Sun May  4 05:21:02 2025

                    Copyright (c) 1991 - 2023 Synopsys, Inc.
   This software and the associated documentation are proprietary to Synopsys,
 Inc. This software may only be used in accordance with the terms and conditions
 of a written license agreement with Synopsys, Inc. All other use, reproduction,
   or distribution of this software is strictly prohibited.  Licensed Products
     communicate with Synopsys servers for the purpose of providing software
    updates, detecting software piracy and verifying that customers are using
    Licensed Products in conformity with the applicable License Key for such
  Licensed Products. Synopsys will use information gathered in connection with
    this process to deliver software updates and pursue software pirates and
                                   infringers.

 Inclusivity & Diversity - Visit SolvNetPlus to read the "Synopsys Statement on
            Inclusivity and Diversity" (Refer to article 000036315 at
                        https://solvnetplus.synopsys.com)

Parsing design file 'design.sv'
Parsing design file 'testbench.sv'
Top Level Modules:
       concurrent_example
TimeScale is 1 ns / 1 ns
Starting vcs inline pass...

1 module and 0 UDP read.
recompiling module concurrent_example
rm -f _cuarc*.so _csrc*.so pre_vcsobj_*.so share_vcsobj_*.so
if [ -x ../simv ]; then chmod a-x ../simv; fi
g++  -o ../simv      -rdynamic  -Wl,-rpath='$ORIGIN'/simv.daidir -Wl,-rpath=./simv.daidir -Wl,-rpath=/apps/vcsmx/vcs/U-2023.03-SP2/linux64/lib -L/apps/vcsmx/vcs/U-2023.03-SP2/linux64/lib  -Wl,-rpath-link=./   objs/amcQw_d.o   _331_archive_1.so   SIM_l.o       rmapats_mop.o rmapats.o rmar.o rmar_nd.o  rmar_llvm_0_1.o rmar_llvm_0_0.o            -lvirsim -lerrorinf -lsnpsmalloc -lvfs    -lvcsnew -lsimprofile -luclinative /apps/vcsmx/vcs/U-2023.03-SP2/linux64/lib/vcs_tls.o   -Wl,-whole-archive  -lvcsucli    -Wl,-no-whole-archive          /apps/vcsmx/vcs/U-2023.03-SP2/linux64/lib/vcs_save_restore_new.o -ldl  -lc -lm -lpthread -ldl 
../simv up to date
CPU time: .471 seconds to compile + .439 seconds to elab + .386 seconds to link
Chronologic VCS simulator copyright 1991-2023
Contains Synopsys proprietary information.
Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  May  4 05:21 2025
PASSED at TIME=5 with a=0 b= 0 
PASSED at TIME=15 with a=1 b= 0 
"testbench.sv", 36: concurrent_example.P1: started at 25ns failed at 25ns
	Offending '(a == b)'
Error: "testbench.sv", 36: concurrent_example.P1: at time 25 ns
FAILED at TIME=25 with a=0 b= 1 
"testbench.sv", 36: concurrent_example.P1: started at 35ns failed at 35ns
	Offending '(a == b)'
Error: "testbench.sv", 36: concurrent_example.P1: at time 35 ns
FAILED at TIME=35 with a=0 b= 1 
"testbench.sv", 36: concurrent_example.P1: started at 45ns failed at 45ns
	Offending '(a == b)'
Error: "testbench.sv", 36: concurrent_example.P1: at time 45 ns
FAILED at TIME=45 with a=0 b= 0 
PASSED at TIME=55 with a=0 b= 1 
"testbench.sv", 36: concurrent_example.P1: started at 65ns failed at 65ns
	Offending '(a == b)'
Error: "testbench.sv", 36: concurrent_example.P1: at time 65 ns
FAILED at TIME=65 with a=0 b= 0 
PASSED at TIME=75 with a=0 b= 0 
PASSED at TIME=85 with a=1 b= 0 
"testbench.sv", 36: concurrent_example.P1: started at 95ns failed at 95ns
	Offending '(a == b)'
Error: "testbench.sv", 36: concurrent_example.P1: at time 95 ns
FAILED at TIME=95 with a=0 b= 1 
"testbench.sv", 36: concurrent_example.P1: started at 105ns failed at 105ns
	Offending '(a == b)'
Error: "testbench.sv", 36: concurrent_example.P1: at time 105 ns
FAILED at TIME=105 with a=0 b= 0 
PASSED at TIME=115 with a=0 b= 1 
"testbench.sv", 36: concurrent_example.P1: started at 125ns failed at 125ns
	Offending '(a == b)'
Error: "testbench.sv", 36: concurrent_example.P1: at time 125 ns
FAILED at TIME=125 with a=0 b= 0 
PASSED at TIME=135 with a=0 b= 1 
"testbench.sv", 36: concurrent_example.P1: started at 145ns failed at 145ns
	Offending '(a == b)'
Error: "testbench.sv", 36: concurrent_example.P1: at time 145 ns
FAILED at TIME=145 with a=0 b= 0 
PASSED at TIME=155 with a=0 b= 0 
$finish called from file "testbench.sv", line 27.
$finish at simulation time                  165
           V C S   S i m u l a t i o n   R e p o r t 
Time: 165 ns
CPU Time:      0.490 seconds;       Data structure size:   0.0Mb
Sun May  4 05:21:04 2025
Finding VCD file...
./waveform.vcd
[2025-05-04 09:21:04 UTC] Opening EPWave...
Done
  
